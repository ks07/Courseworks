module encrypt_v3( input  wire            clk,

                   input  wire [ 79 : 0 ]   K,
                   input  wire [ 63 : 0 ]   M,
                   output wire [ 63 : 0 ]   C );

  // fill in this module with solution

endmodule
