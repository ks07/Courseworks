module round( output wire [ 63 : 0 ] r, 
              input  wire [ 63 : 0 ] x, 
              input  wire [ 79 : 0 ] k );

  // fill in this module with solution

endmodule
