module encrypt_v2( input  wire            clk,
                   input  wire            req,
                   output wire            ack,

                   input  wire [ 79 : 0 ]   K,
                   input  wire [ 63 : 0 ]   M,
                   output wire [ 63 : 0 ]   C );

  // fill in this module with solution

endmodule
