module key_schedule( output wire [ 79 : 0 ] r,
                     input  wire [ 79 : 0 ] x,
                     input  wire [  4 : 0 ] i );

  // fill in this module with solution

endmodule
