module encrypt_v1( input  wire [ 79 : 0 ]   K,
                   input  wire [ 63 : 0 ]   M,
                   output wire [ 63 : 0 ]   C );

  // fill in this module with solution

endmodule
