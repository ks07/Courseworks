library verilog;
use verilog.vl_types.all;
entity calc1_reference_test is
end calc1_reference_test;
