module clr_28bit( output wire [ 27 : 0 ] r,
                  input  wire [ 27 : 0 ] x,
                  input  wire [  3 : 0 ] y );

  // fill in this module with solution

endmodule
