module sbox( output wire [ 3 : 0 ] r,
             input  wire [ 3 : 0 ] x );

  // fill in this module with solution

endmodule                
